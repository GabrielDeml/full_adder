module halfAdder(
    input 
)